---------------------------------------------------------------------------
--
--  File        : buf_bsram.vhd
--
--  Title       : BSRAM for configurable size data buffer
--
--  Author      : Jukka Pietarinen
--                Micro-Research Finland Oy
--                <jukka.pietarinen@mrf.fi>
--
--  Description :
--
---------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
-- LIBRARY UNISIM;
-- use UNISIM.VCOMPONENTS.ALL;

entity buf_bsram IS
  port (
    addra: IN std_logic_VECTOR(10 downto 0);
    addrb: IN std_logic_VECTOR(8 downto 0);
    clka: IN std_logic;
    clkb: IN std_logic;
    dina: IN std_logic_VECTOR(7 downto 0);
    doutb: OUT std_logic_VECTOR(31 downto 0);
    wea: IN std_logic);
end buf_bsram;

architecture structure of buf_bsram is

  signal vcc : std_logic;
  signal gnd : std_logic;
  signal gnd8 : std_logic_vector(7 downto 0);
  signal gnd32 : std_logic_vector(31 downto 0);

  signal douta: std_logic_VECTOR(7 downto 0);
  signal dinb: std_logic_VECTOR(31 downto 0) := (others => '0');
  signal web: std_logic := '0';
  
  component RAMB16_S9_S36 is
    generic (
      INIT_00 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_A : bit_vector  := X"000";
      INIT_B : bit_vector  := X"000";
      INITP_00 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_01 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_02 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_03 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_04 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_05 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_06 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_07 : bit_vector :=
      X"0000000000000000000000000000000000000000000000000000000000000000";
      SRVAL_A : bit_vector  := X"000";
      SRVAL_B : bit_vector  := X"000";
      WRITE_MODE_A : string := "WRITE_FIRST";
      WRITE_MODE_B : string := "WRITE_FIRST"
      );

    port (
      DOA   : out std_logic_vector(7 downto 0);
      DOB   : out std_logic_vector(31 downto 0);
      DOPA  : out std_logic_vector(0 downto 0);
      DOPB  : out std_logic_vector(3 downto 0);
      ADDRA : in  std_logic_vector(10 downto 0);
      ADDRB : in  std_logic_vector(8 downto 0);
      CLKA  : in  std_ulogic;
      CLKB  : in  std_ulogic;
      DIA   : in  std_logic_vector(7 downto 0);
      DIB   : in  std_logic_vector(31 downto 0);
      DIPA  : in  std_logic_vector(0 downto 0);
      DIPB  : in  std_logic_vector(3 downto 0);
      ENA   : in  std_ulogic;
      ENB   : in  std_ulogic;
      SSRA  : in  std_ulogic;
      SSRB  : in  std_ulogic;
      WEA   : in  std_ulogic;
      WEB   : in  std_ulogic);
  end component;
  
begin

  vcc <= '1';
  gnd <= '0';
  gnd8 <= (others => '0');
  gnd32 <= (others => '0');

  i_bsram : RAMB16_S9_S36
    port map (
      DOA => douta,
      DOB => doutb,
      DOPA => open,
      DOPB => open,
      ADDRA => addra,
      ADDRB => addrb,
      CLKA => clka,
      CLKB => clkb,
      DIA => dina,
      DIB => dinb,
      DIPA => gnd8(0 downto 0),
      DIPB => gnd8(3 downto 0),
      ENA => vcc,
      ENB => vcc,
      SSRA => gnd,
      SSRB => gnd,
      WEA => wea,
      WEB => web);

end structure;
